"0111100110011100000000111111101111111111111111111111111000111111000111111000011111110001100100000000" &
"1110001101001001111100111111001000000000000000000000101000001000000100001110111111111011110111101001" &
"0111111111111100011111000000111100000011011110001110011101100011111000111111100000111001110000110110" &
"1011100011000011111110011111110111000101111110001111110011111110011110111101110001111110001111100000" &
"1111000011101001000100011110000001010000000010000000001000000000110000000011100000001111110000111110" &
"1110111110101011111100001011110000011111000000111110000000011011100000111100000011111000001111110001" &
"1111101000011111100011111100001111000000111010000111100101111110001110100000111110100111111000110100" &
"0010011111111111111101110010110100000000000110000000001000010000001100000111110100111111011111111101" &

"0111111111100111111101111101110001111111000011111100111111010011110000000010000110111101000111011000" &
"0010100101111011110011110001111001100111101000011111110000101100000101100000001110000110110011000011" &
"0111110100111111111110111111111110010111011000001111100001100110011100111001111011000110010011100000" &
"0011111111000011111100110101101011100001000110011010111100010000000000000110001110110011100001000101" &
"0000000001010000000011100000010110000001111100011011010001101101000110000010110110010001100000000010" &
"1110100000111100000001110000001000100001000000010000000000000000100010000000011100001111010000011110" &
"1000000011000110111100110000000010000000000100000000110000000001100110011110011111111000011111100011" &
"0000000000110000000011000000001110010000111010000011000100011110010011111010010010000010100000001000" &

"1001011111000000101100001011110000011111000000101000000110001111000000111100000011111000001010000000" &
"1101110011101101011011100010001100000000111001111001101111111101110111010111011100011110001101111011" &
"1100001110000000111101100001111000011111101111111111111011111111110000111110000010011000000011100000" &
"1110001110111001111110000011010000000111000001100000001111001100111000110011110000000111001000001110" &
"1110101111111111111111111100011111000001111110000011111101111111011111000101111100001111100011111110" &
"0111111110001111111000011111100000100101001111000000010000000001001000001111110101111111110111111110" &
"1111100000010010000000000000000010000000011111110111111111111111011101111110111111110001111110000000" &
"1111111100011110110010011010001111110000111111001011111100000001110111000001111100010111110011111111" &

"0000010111100001111100000011110100000011010100100000000100010000000111000001111100000011110000100111" &
"0001111111000000101110000000001100001111010001111010111010010110101011010011000010001001111100011111" &
"1000001110000001111100000111110000111111000100110111111010111111111111111111111101111111110011111111" &
"0010111011111001111110000011110000001111010111100000000011010000101111000001111110000110110000000010" &
"1111111111111110000101110000011111000011111110011111111111111111000101111100000111111000010011111111" &
"0011111111011111111000111111110000111111000001111000011111001100101111110000111110001011011000000100" &
"1110100000110111101000001111110001111111000111011100111111100000000100000000111100001111100011111111" &
"1101101000111111000011111110001111111110100011111010001111111111111110111111100011111110001111111000" &

"0011110110111111111111111111110111111111111000010100000001000000001010000001000101011111000001101111" &
"1100010001010011011011111111101011111111001111111010111011110110001110110100000000000011100001000011" &
"0111111111111111111111111111110111111111111111101100000000110000000001000000001101100110011110000000" &
"1011111111111111111100111111101111111100111110011011001111011000000000000100000000100011110011101110" &
"1000100001000000000000000000000000100001000111000100001000010011000101000101001101100000011010100000" &
"1000000000110000000011000000001110100000110111100011111011000110111010000011110000010011001000001100" &
"0000000001000000001100001111111111011011111001101111101111111100110010011010000011101000000111000000" &
"0100000001000000000010000000000000000000100100100000110010110110010011011100010111000000101010000111" &

"1111010000111100000011110000001100000000110110000000000100100000000111000000011100000111111000000011" &
"1111111011111111111101110000011000000000111010000011111010111100001011110000000111000111101110001111" &
"0011110011111100000010110000001101000000011000000011101001111110111111011111111100111111110001111110" &
"1011000000010000000101100000001111000000001111100000011001110000001111100001111110000000101000000011" &
"1101111111100011111010001111111000011111100011111111001111111111011100111111001011111000001100111110" &
"0100000000110000001110110000001011110001111100110011111111101111111111110010110011011000000001000000" &
"0000111111010011111111100000011111001000101000000000010000000000000000000111001100011111110011011110" &
"0000011111000011111100001111110000001111000010111111111100000111111000111111100011111110001111110000" &

"1111111111111111100011111000001111100001111110000111110110111111111011111101111111111111101010000010" &
"0000000000001000000000011111100011111110101111111000111111000000011100010100010110000010001101100000" &
"0111111000011111100111111111111111111011011111101101011111000000110100000111100110000001111000000010" &
"1011111000001110000001111000001111100001011011011111111111111111001110111101111001111110010000000000" &
"0000000000000000111000000011100000011111000001111100000111000000101100100011111111000111011100011110" &
"1000000111000000000100000000000000000011000000001110001111111111111110011111110101111111001001110011" &
"1110111111101101110000100001101110001100101100001011111111101111010110011111111100000011100000011101" &
"0000000010000001111100001111110000001111000000111100001010110000011101000110110100111110000111111110" &

"0000000000000000001000000000010000000001000110100100010001100011110111111111011111111111011111111001" &
"1001111011111011011010111111110110000110110000011110001100011001110011111100001011100011110101110000" &
"1111111100000000111100000001110000000011000000001100011000100111100001111110001111110110111111111111" &
"1000000010100000000111100011111000000001100000010010000111011000011111000011111101011000001011101111" &
"0011111011011111111001001101011111101011010110011100011000010011010001001101001111000001111110000011" &
"1100000100111111000011001110101000111011000001110000000100100000000000000010000000000000000000000000" &
"0000011001100001101110000000110000000000110101101000011101111011111111000011110000111000001111110001" &
"1111111111010111101011110010011111000000110100100011000001111110000111111000000011100000100000000000" &

"1111111010001011110000110001100111001111111110100001011110001111111111111110111111110011111111111110" &
"0000100000001001011001011100000010001110011111111010111111100011011100001111110010010100000011111100" &
"0011101111001111111110111110011100011111100001111000100110001100111001111101111111011111110000001111" &
"0000001100010111111001110010111111101101001101111000111100000011110000111100111101111111111111111010" &
"1001111011001111111001101110101010011100110001111011000111110000111110000100100000000110001000111000" &
"0000011110001111111111111111111111101111111111111110101101000010111101000111110101111111111111111110" &
"1010111101011110101001110011011100001111100001111100011111101111100000111110000111100111110000111111" &
"0011111101101011111100001111110000111101011110111011111111111100101111000001100100001100000001110111" &

"0111000000011101100011111111011111111011111010111111000111111100011110100101111100101111101000111110" &
"1100100000000100000000110000000011000000011111000001111101011011110000100011111000000001000100010100" &
"0011101000011100111111100001111110111111100000011100000010110000001111000000011110110010111110111110" &
"0100001110010011111111111101111111101111111111101110011000000011000001010101001000000000001000001111" &
"0110111110111111111111111111100011110010000111100100011100011111100000111100001011110000001101110000" &
"0001010101000111111100001111110011111110111001111111110101001111011000111001100001100111000000000011" &
"1111111000011111100011111000001111111101100001010010001011000000011000000011100000001000011111110001" &
"1111111011111111111110111111110000011000000101000001010100101111100010111100000011100000000000000100" &

