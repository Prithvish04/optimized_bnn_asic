"000000000" &
"100010000" &
"001111010" &
"111111111" &
"111111111" &
"011111111" &
"000000001" &
"000100100" &
"010000010" &

"000000000" &
"000010000" &
"000100100" &
"111001110" &
"011001100" &
"111110001" &
"011010010" &
"001000001" &
"000000100" &

"111110000" &
"001000000" &
"000000000" &
"000000000" &
"000000000" &
"100110000" &
"111111111" &
"111111111" &
"111111110" &

"000000010" &
"010000000" &
"000001100" &
"000111111" &
"101111111" &
"111111111" &
"111111101" &
"101000010" &
"000000000" &

"110000000" &
"011000011" &
"111000101" &
"111010001" &
"011000011" &
"111000001" &
"011010011" &
"011100011" &
"000000110" &

"111110011" &
"111110001" &
"110111100" &
"000111100" &
"001111100" &
"111011111" &
"100001111" &
"100010111" &
"001110011" &

"111100011" &
"101000011" &
"110001111" &
"100011111" &
"000111110" &
"001111110" &
"111111100" &
"111110011" &
"111000101" &

"010001100" &
"100011100" &
"001111010" &
"010011100" &
"000111000" &
"011111010" &
"000111000" &
"001111010" &
"010111100" &

