"0000000000000000000000000000" &
"0000000000000000000000000000" &
"0000000000000000000000000000" &
"0000000000000000000000000000" &
"0000000000001111100000000000" &
"0000000000111111110000000000" &
"0000000001111111110000000000" &
"0000000000000001110000000000" &
"0000000000000011110000000000" &
"0000000000000011100000000000" &
"0000000000000111000000000000" &
"0000000000001110000000000000" &
"0000000000011111000000000000" &
"0000000000011111100000000000" &
"0000000000000111110000000000" &
"0000000000000001111000000000" &
"0000000000000000111000000000" &
"0000000000000000011100000000" &
"0000000000000000011100000000" &
"0000000000000000011100000000" &
"0000000011000001111000000000" &
"0000000011111111110000000000" &
"0000000011111111100000000000" &
"0000000000111000000000000000" &
"0000000000000000000000000000" &
"0000000000000000000000000000" &
"0000000000000000000000000000" &
"0000000000000000000000000000" &
