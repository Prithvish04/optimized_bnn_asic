	px_0: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(0));
	px_1: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(1));
	px_2: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(2));
	px_3: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(3));
	px_4: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(4));
	px_5: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(5));
	px_6: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(6));
	px_7: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(7));
	px_8: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(8));
	px_9: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(9));
	px_10: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(10));
	px_11: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(11));
	px_12: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(12));
	px_13: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(13));
	px_14: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(14));
	px_15: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(15));
	px_16: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(16));
	px_17: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(17));
	px_18: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(18));
	px_19: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(19));
	px_20: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(20));
	px_21: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(21));
	px_22: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(22));
	px_23: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(23));
	px_24: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(24));
	px_25: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(25));
	px_26: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(26));
	px_27: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(27));
	px_28: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(28));
	px_29: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(29));
	px_30: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(30));
	px_31: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(31));
	px_32: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(32));
	px_33: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(33));
	px_34: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(34));
	px_35: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(35));
	px_36: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(36));
	px_37: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(37));
	px_38: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(38));
	px_39: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(39));
	px_40: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(40));
	px_41: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(41));
	px_42: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(42));
	px_43: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(43));
	px_44: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(44));
	px_45: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(45));
	px_46: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(46));
	px_47: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(47));
	px_48: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(48));
	px_49: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(49));
	px_50: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(50));
	px_51: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(51));
	px_52: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(52));
	px_53: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(53));
	px_54: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(54));
	px_55: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(55));
	px_56: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(56));
	px_57: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(57));
	px_58: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(58));
	px_59: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(59));
	px_60: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(60));
	px_61: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(61));
	px_62: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(62));
	px_63: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(63));
	px_64: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(64));
	px_65: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(65));
	px_66: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(66));
	px_67: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(67));
	px_68: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(68));
	px_69: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(69));
	px_70: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(70));
	px_71: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(71));
	px_72: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(72));
	px_73: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(73));
	px_74: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(74));
	px_75: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(75));
	px_76: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(76));
	px_77: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(77));
	px_78: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(78));
	px_79: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(79));
	px_80: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(80));
	px_81: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(81));
	px_82: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(82));
	px_83: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(83));
	px_84: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(84));
	px_85: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(85));
	px_86: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(86));
	px_87: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(87));
	px_88: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(88));
	px_89: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(89));
	px_90: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(90));
	px_91: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(91));
	px_92: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(92));
	px_93: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(93));
	px_94: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(94));
	px_95: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(95));
	px_96: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(96));
	px_97: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(97));
	px_98: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(98));
	px_99: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(99));
	px_100: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(100));
	px_101: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(101));
	px_102: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(102));
	px_103: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(103));
	px_104: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(104));
	px_105: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(105));
	px_106: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(106));
	px_107: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(107));
	px_108: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(108));
	px_109: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(109));
	px_110: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(110));
	px_111: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(111));
	px_112: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(112));
	px_113: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(113));
	px_114: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(114));
	px_115: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(115));
	px_116: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(116));
	px_117: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(117));
	px_118: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(118));
	px_119: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(119));
	px_120: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(120));
	px_121: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(121));
	px_122: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(122));
	px_123: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(123));
	px_124: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(124));
	px_125: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(125));
	px_126: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(126));
	px_127: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(127));
	px_128: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(128));
	px_129: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(129));
	px_130: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(130));
	px_131: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(131));
	px_132: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(132));
	px_133: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(133));
	px_134: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(134));
	px_135: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(135));
	px_136: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(136));
	px_137: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(137));
	px_138: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(138));
	px_139: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(139));
	px_140: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(140));
	px_141: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(141));
	px_142: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(142));
	px_143: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(143));
	px_144: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(144));
	px_145: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(145));
	px_146: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(146));
	px_147: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(147));
	px_148: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(148));
	px_149: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(149));
	px_150: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(150));
	px_151: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(151));
	px_152: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(152));
	px_153: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(153));
	px_154: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(154));
	px_155: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(155));
	px_156: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(156));
	px_157: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(157));
	px_158: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(158));
	px_159: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(159));
	px_160: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(160));
	px_161: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(161));
	px_162: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(162));
	px_163: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(163));
	px_164: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(164));
	px_165: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(165));
	px_166: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(166));
	px_167: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(167));
	px_168: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(168));
	px_169: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(169));
	px_170: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(170));
	px_171: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(171));
	px_172: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(172));
	px_173: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(173));
	px_174: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(174));
	px_175: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(175));
	px_176: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(176));
	px_177: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(177));
	px_178: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(178));
	px_179: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(179));
	px_180: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(180));
	px_181: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(181));
	px_182: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(182));
	px_183: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(183));
	px_184: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(184));
	px_185: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(185));
	px_186: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(186));
	px_187: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(187));
	px_188: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(188));
	px_189: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(189));
	px_190: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(190));
	px_191: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(191));
	px_192: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(192));
	px_193: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(193));
	px_194: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(194));
	px_195: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(195));
	px_196: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(196));
	px_197: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(197));
	px_198: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(198));
	px_199: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(199));
	px_200: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(200));
	px_201: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(201));
	px_202: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(202));
	px_203: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(203));
	px_204: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(204));
	px_205: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(205));
	px_206: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(206));
	px_207: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(207));
	px_208: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(208));
	px_209: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(209));
	px_210: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(210));
	px_211: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(211));
	px_212: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(212));
	px_213: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(213));
	px_214: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(214));
	px_215: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(215));
	px_216: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(216));
	px_217: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(217));
	px_218: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(218));
	px_219: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(219));
	px_220: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(220));
	px_221: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(221));
	px_222: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(222));
	px_223: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(223));
	px_224: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(224));
	px_225: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(225));
	px_226: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(226));
	px_227: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(227));
	px_228: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(228));
	px_229: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(229));
	px_230: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(230));
	px_231: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(231));
	px_232: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(232));
	px_233: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(233));
	px_234: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(234));
	px_235: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(235));
	px_236: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(236));
	px_237: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(237));
	px_238: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(238));
	px_239: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(239));
	px_240: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(240));
	px_241: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(241));
	px_242: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(242));
	px_243: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(243));
	px_244: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(244));
	px_245: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(245));
	px_246: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(246));
	px_247: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(247));
	px_248: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(248));
	px_249: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(249));
	px_250: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(250));
	px_251: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(251));
	px_252: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(252));
	px_253: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(253));
	px_254: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(254));
	px_255: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(255));
	px_256: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(256));
	px_257: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(257));
	px_258: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(258));
	px_259: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(259));
	px_260: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(260));
	px_261: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(261));
	px_262: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(262));
	px_263: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(263));
	px_264: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(264));
	px_265: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(265));
	px_266: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(266));
	px_267: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(267));
	px_268: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(268));
	px_269: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(269));
	px_270: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(270));
	px_271: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(271));
	px_272: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(272));
	px_273: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(273));
	px_274: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(274));
	px_275: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(275));
	px_276: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(276));
	px_277: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(277));
	px_278: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(278));
	px_279: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(279));
	px_280: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(280));
	px_281: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(281));
	px_282: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(282));
	px_283: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(283));
	px_284: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(284));
	px_285: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(285));
	px_286: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(286));
	px_287: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(287));
	px_288: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(288));
	px_289: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(289));
	px_290: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(290));
	px_291: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(291));
	px_292: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(292));
	px_293: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(293));
	px_294: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(294));
	px_295: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(295));
	px_296: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(296));
	px_297: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(297));
	px_298: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(298));
	px_299: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(299));
	px_300: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(300));
	px_301: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(301));
	px_302: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(302));
	px_303: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(303));
	px_304: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(304));
	px_305: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(305));
	px_306: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(306));
	px_307: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(307));
	px_308: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(308));
	px_309: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(309));
	px_310: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(310));
	px_311: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(311));
	px_312: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(312));
	px_313: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(313));
	px_314: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(314));
	px_315: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(315));
	px_316: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(316));
	px_317: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(317));
	px_318: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(318));
	px_319: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(319));
	px_320: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(320));
	px_321: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(321));
	px_322: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(322));
	px_323: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(323));
	px_324: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(324));
	px_325: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(325));
	px_326: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(326));
	px_327: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(327));
	px_328: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(328));
	px_329: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(329));
	px_330: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(330));
	px_331: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(331));
	px_332: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(332));
	px_333: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(333));
	px_334: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(334));
	px_335: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(335));
	px_336: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(336));
	px_337: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(337));
	px_338: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(338));
	px_339: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(339));
	px_340: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(340));
	px_341: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(341));
	px_342: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(342));
	px_343: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(343));
	px_344: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(344));
	px_345: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(345));
	px_346: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(346));
	px_347: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(347));
	px_348: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(348));
	px_349: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(349));
	px_350: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(350));
	px_351: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(351));
	px_352: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(352));
	px_353: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(353));
	px_354: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(354));
	px_355: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(355));
	px_356: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(356));
	px_357: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(357));
	px_358: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(358));
	px_359: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(359));
	px_360: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(360));
	px_361: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(361));
	px_362: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(362));
	px_363: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(363));
	px_364: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(364));
	px_365: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(365));
	px_366: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(366));
	px_367: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(367));
	px_368: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(368));
	px_369: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(369));
	px_370: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(370));
	px_371: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(371));
	px_372: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(372));
	px_373: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(373));
	px_374: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(374));
	px_375: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(375));
	px_376: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(376));
	px_377: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(377));
	px_378: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(378));
	px_379: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(379));
	px_380: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(380));
	px_381: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(381));
	px_382: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(382));
	px_383: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(383));
	px_384: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(384));
	px_385: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(385));
	px_386: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(386));
	px_387: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(387));
	px_388: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(388));
	px_389: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(389));
	px_390: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(390));
	px_391: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(391));
	px_392: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(392));
	px_393: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(393));
	px_394: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(394));
	px_395: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(395));
	px_396: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(396));
	px_397: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(397));
	px_398: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(398));
	px_399: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(399));
	px_400: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(400));
	px_401: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(401));
	px_402: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(402));
	px_403: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(403));
	px_404: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(404));
	px_405: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(405));
	px_406: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(406));
	px_407: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(407));
	px_408: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(408));
	px_409: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(409));
	px_410: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(410));
	px_411: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(411));
	px_412: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(412));
	px_413: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(413));
	px_414: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(414));
	px_415: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(415));
	px_416: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(416));
	px_417: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(417));
	px_418: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(418));
	px_419: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(419));
	px_420: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(420));
	px_421: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(421));
	px_422: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(422));
	px_423: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(423));
	px_424: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(424));
	px_425: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(425));
	px_426: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(426));
	px_427: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(427));
	px_428: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(428));
	px_429: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(429));
	px_430: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(430));
	px_431: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(431));
	px_432: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(432));
	px_433: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(433));
	px_434: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(434));
	px_435: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(435));
	px_436: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(436));
	px_437: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(437));
	px_438: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(438));
	px_439: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(439));
	px_440: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(440));
	px_441: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(441));
	px_442: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(442));
	px_443: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(443));
	px_444: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(444));
	px_445: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(445));
	px_446: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(446));
	px_447: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(447));
	px_448: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(448));
	px_449: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(449));
	px_450: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(450));
	px_451: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(451));
	px_452: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(452));
	px_453: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(453));
	px_454: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(454));
	px_455: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(455));
	px_456: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(456));
	px_457: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(457));
	px_458: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(458));
	px_459: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(459));
	px_460: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(460));
	px_461: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(461));
	px_462: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(462));
	px_463: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(463));
	px_464: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(464));
	px_465: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(465));
	px_466: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(466));
	px_467: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(467));
	px_468: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(468));
	px_469: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(469));
	px_470: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(470));
	px_471: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(471));
	px_472: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(472));
	px_473: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(473));
	px_474: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(474));
	px_475: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(475));
	px_476: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(476));
	px_477: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(477));
	px_478: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(478));
	px_479: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(479));
	px_480: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(480));
	px_481: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(481));
	px_482: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(482));
	px_483: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(483));
	px_484: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(484));
	px_485: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(485));
	px_486: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(486));
	px_487: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(487));
	px_488: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(488));
	px_489: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(489));
	px_490: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(490));
	px_491: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(491));
	px_492: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(492));
	px_493: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(493));
	px_494: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(494));
	px_495: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(495));
	px_496: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(496));
	px_497: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(497));
	px_498: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(498));
	px_499: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(499));
	px_500: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(500));
	px_501: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(501));
	px_502: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(502));
	px_503: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(503));
	px_504: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(504));
	px_505: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(505));
	px_506: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(506));
	px_507: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(507));
	px_508: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(508));
	px_509: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(509));
	px_510: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(510));
	px_511: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(511));
	px_512: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(512));
	px_513: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(513));
	px_514: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(514));
	px_515: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(515));
	px_516: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(516));
	px_517: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(517));
	px_518: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(518));
	px_519: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(519));
	px_520: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(520));
	px_521: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(521));
	px_522: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(522));
	px_523: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(523));
	px_524: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(524));
	px_525: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(525));
	px_526: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(526));
	px_527: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(527));
	px_528: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(528));
	px_529: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(529));
	px_530: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(530));
	px_531: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(531));
	px_532: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(532));
	px_533: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(533));
	px_534: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(534));
	px_535: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(535));
	px_536: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(536));
	px_537: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(537));
	px_538: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(538));
	px_539: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(539));
	px_540: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(540));
	px_541: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(541));
	px_542: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(542));
	px_543: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(543));
	px_544: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(544));
	px_545: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(545));
	px_546: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(546));
	px_547: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(547));
	px_548: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(548));
	px_549: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(549));
	px_550: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(550));
	px_551: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(551));
	px_552: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(552));
	px_553: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(553));
	px_554: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(554));
	px_555: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(555));
	px_556: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(556));
	px_557: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(557));
	px_558: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(558));
	px_559: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(559));
	px_560: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(560));
	px_561: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(561));
	px_562: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(562));
	px_563: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(563));
	px_564: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(564));
	px_565: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(565));
	px_566: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(566));
	px_567: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(567));
	px_568: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(568));
	px_569: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(569));
	px_570: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(570));
	px_571: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(571));
	px_572: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(572));
	px_573: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(573));
	px_574: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(574));
	px_575: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(575));
	px_576: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(576));
	px_577: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(577));
	px_578: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(578));
	px_579: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(579));
	px_580: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(580));
	px_581: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(581));
	px_582: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(582));
	px_583: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(583));
	px_584: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(584));
	px_585: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(585));
	px_586: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(586));
	px_587: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(587));
	px_588: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(588));
	px_589: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(589));
	px_590: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(590));
	px_591: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(591));
	px_592: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(592));
	px_593: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(593));
	px_594: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(594));
	px_595: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(595));
	px_596: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(596));
	px_597: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(597));
	px_598: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(598));
	px_599: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(599));
	px_600: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(600));
	px_601: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(601));
	px_602: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(602));
	px_603: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(603));
	px_604: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(604));
	px_605: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(605));
	px_606: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(606));
	px_607: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(607));
	px_608: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(608));
	px_609: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(609));
	px_610: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(610));
	px_611: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(611));
	px_612: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(612));
	px_613: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(613));
	px_614: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(614));
	px_615: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(615));
	px_616: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(616));
	px_617: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(617));
	px_618: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(618));
	px_619: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(619));
	px_620: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(620));
	px_621: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(621));
	px_622: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(622));
	px_623: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(623));
	px_624: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(624));
	px_625: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(625));
	px_626: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(626));
	px_627: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(627));
	px_628: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(628));
	px_629: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(629));
	px_630: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(630));
	px_631: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(631));
	px_632: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(632));
	px_633: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(633));
	px_634: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(634));
	px_635: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(635));
	px_636: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(636));
	px_637: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(637));
	px_638: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(638));
	px_639: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(639));
	px_640: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(640));
	px_641: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(641));
	px_642: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(642));
	px_643: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(643));
	px_644: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(644));
	px_645: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(645));
	px_646: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(646));
	px_647: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(647));
	px_648: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(648));
	px_649: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(649));
	px_650: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(650));
	px_651: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(651));
	px_652: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(652));
	px_653: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(653));
	px_654: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(654));
	px_655: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(655));
	px_656: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_px(656));
	px_657: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(657));
	px_658: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(658));
	px_659: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(659));
	px_660: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(660));
	px_661: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(661));
	px_662: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(662));
	px_663: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(663));
	px_664: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(664));
	px_665: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(665));
	px_666: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(666));
	px_667: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(667));
	px_668: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(668));
	px_669: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(669));
	px_670: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(670));
	px_671: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(671));
	px_672: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(672));
	px_673: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(673));
	px_674: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(674));
	px_675: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(675));
	px_676: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(676));
	px_677: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(677));
	px_678: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(678));
	px_679: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(679));
	px_680: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(680));
	px_681: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(681));
	px_682: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(682));
	px_683: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(683));
	px_684: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(684));
	px_685: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(685));
	px_686: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(686));
	px_687: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(687));
	px_688: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(688));
	px_689: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(689));
	px_690: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(690));
	px_691: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(691));
	px_692: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(692));
	px_693: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(693));
	px_694: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(694));
	px_695: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(695));
	px_696: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(696));
	px_697: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(697));
	px_698: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(698));
	px_699: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(699));
	px_700: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(700));
	px_701: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(701));
	px_702: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(702));
	px_703: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(703));
	px_704: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(704));
	px_705: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(705));
	px_706: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(706));
	px_707: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(707));
	px_708: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(708));
	px_709: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(709));
	px_710: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(710));
	px_711: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(711));
	px_712: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(712));
	px_713: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(713));
	px_714: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(714));
	px_715: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(715));
	px_716: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(716));
	px_717: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(717));
	px_718: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(718));
	px_719: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(719));
	px_720: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(720));
	px_721: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(721));
	px_722: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(722));
	px_723: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(723));
	px_724: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(724));
	px_725: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(725));
	px_726: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(726));
	px_727: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(727));
	px_728: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(728));
	px_729: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(729));
	px_730: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(730));
	px_731: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(731));
	px_732: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(732));
	px_733: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(733));
	px_734: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(734));
	px_735: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(735));
	px_736: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(736));
	px_737: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(737));
	px_738: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(738));
	px_739: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(739));
	px_740: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(740));
	px_741: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(741));
	px_742: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(742));
	px_743: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(743));
	px_744: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(744));
	px_745: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(745));
	px_746: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(746));
	px_747: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(747));
	px_748: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(748));
	px_749: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(749));
	px_750: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(750));
	px_751: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(751));
	px_752: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(752));
	px_753: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(753));
	px_754: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(754));
	px_755: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(755));
	px_756: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(756));
	px_757: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(757));
	px_758: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(758));
	px_759: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(759));
	px_760: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(760));
	px_761: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(761));
	px_762: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(762));
	px_763: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(763));
	px_764: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(764));
	px_765: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(765));
	px_766: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(766));
	px_767: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(767));
	px_768: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(768));
	px_769: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(769));
	px_770: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(770));
	px_771: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(771));
	px_772: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(772));
	px_773: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(773));
	px_774: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(774));
	px_775: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(775));
	px_776: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(776));
	px_777: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(777));
	px_778: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(778));
	px_779: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(779));
	px_780: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(780));
	px_781: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(781));
	px_782: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(782));
	px_783: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_px(783));
