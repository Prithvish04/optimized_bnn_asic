	conv_row_0: 	reg_8bit port map (CLK => CLK, rst => '0', input => "000000000", output => elem_conv_row(0));
	conv_row_1: 	reg_8bit port map (CLK => CLK, rst => '0', input => "100010000", output => elem_conv_row(1));
	conv_row_2: 	reg_8bit port map (CLK => CLK, rst => '0', input => "001111010", output => elem_conv_row(2));
	conv_row_3: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111111111", output => elem_conv_row(3));
	conv_row_4: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111111111", output => elem_conv_row(4));
	conv_row_5: 	reg_8bit port map (CLK => CLK, rst => '0', input => "011111111", output => elem_conv_row(5));
	conv_row_6: 	reg_8bit port map (CLK => CLK, rst => '0', input => "000000001", output => elem_conv_row(6));
	conv_row_7: 	reg_8bit port map (CLK => CLK, rst => '0', input => "000100100", output => elem_conv_row(7));
	conv_row_8: 	reg_8bit port map (CLK => CLK, rst => '0', input => "010000010", output => elem_conv_row(8));

	conv_row_9: 	reg_8bit port map (CLK => CLK, rst => '0', input => "000000000", output => elem_conv_row(9));
	conv_row_10: 	reg_8bit port map (CLK => CLK, rst => '0', input => "000010000", output => elem_conv_row(10));
	conv_row_11: 	reg_8bit port map (CLK => CLK, rst => '0', input => "000100100", output => elem_conv_row(11));
	conv_row_12: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111001110", output => elem_conv_row(12));
	conv_row_13: 	reg_8bit port map (CLK => CLK, rst => '0', input => "011001100", output => elem_conv_row(13));
	conv_row_14: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111110001", output => elem_conv_row(14));
	conv_row_15: 	reg_8bit port map (CLK => CLK, rst => '0', input => "011010010", output => elem_conv_row(15));
	conv_row_16: 	reg_8bit port map (CLK => CLK, rst => '0', input => "001000001", output => elem_conv_row(16));
	conv_row_17: 	reg_8bit port map (CLK => CLK, rst => '0', input => "000000100", output => elem_conv_row(17));

	conv_row_18: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111110000", output => elem_conv_row(18));
	conv_row_19: 	reg_8bit port map (CLK => CLK, rst => '0', input => "001000000", output => elem_conv_row(19));
	conv_row_20: 	reg_8bit port map (CLK => CLK, rst => '0', input => "000000000", output => elem_conv_row(20));
	conv_row_21: 	reg_8bit port map (CLK => CLK, rst => '0', input => "000000000", output => elem_conv_row(21));
	conv_row_22: 	reg_8bit port map (CLK => CLK, rst => '0', input => "000000000", output => elem_conv_row(22));
	conv_row_23: 	reg_8bit port map (CLK => CLK, rst => '0', input => "100110000", output => elem_conv_row(23));
	conv_row_24: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111111111", output => elem_conv_row(24));
	conv_row_25: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111111111", output => elem_conv_row(25));
	conv_row_26: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111111110", output => elem_conv_row(26));

	conv_row_27: 	reg_8bit port map (CLK => CLK, rst => '0', input => "000000010", output => elem_conv_row(27));
	conv_row_28: 	reg_8bit port map (CLK => CLK, rst => '0', input => "010000000", output => elem_conv_row(28));
	conv_row_29: 	reg_8bit port map (CLK => CLK, rst => '0', input => "000001100", output => elem_conv_row(29));
	conv_row_30: 	reg_8bit port map (CLK => CLK, rst => '0', input => "000111111", output => elem_conv_row(30));
	conv_row_31: 	reg_8bit port map (CLK => CLK, rst => '0', input => "101111111", output => elem_conv_row(31));
	conv_row_32: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111111111", output => elem_conv_row(32));
	conv_row_33: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111111101", output => elem_conv_row(33));
	conv_row_34: 	reg_8bit port map (CLK => CLK, rst => '0', input => "101000010", output => elem_conv_row(34));
	conv_row_35: 	reg_8bit port map (CLK => CLK, rst => '0', input => "000000000", output => elem_conv_row(35));

	conv_row_36: 	reg_8bit port map (CLK => CLK, rst => '0', input => "110000000", output => elem_conv_row(36));
	conv_row_37: 	reg_8bit port map (CLK => CLK, rst => '0', input => "011000011", output => elem_conv_row(37));
	conv_row_38: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111000101", output => elem_conv_row(38));
	conv_row_39: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111010001", output => elem_conv_row(39));
	conv_row_40: 	reg_8bit port map (CLK => CLK, rst => '0', input => "011000011", output => elem_conv_row(40));
	conv_row_41: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111000001", output => elem_conv_row(41));
	conv_row_42: 	reg_8bit port map (CLK => CLK, rst => '0', input => "011010011", output => elem_conv_row(42));
	conv_row_43: 	reg_8bit port map (CLK => CLK, rst => '0', input => "011100011", output => elem_conv_row(43));
	conv_row_44: 	reg_8bit port map (CLK => CLK, rst => '0', input => "000000110", output => elem_conv_row(44));

	conv_row_45: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111110011", output => elem_conv_row(45));
	conv_row_46: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111110001", output => elem_conv_row(46));
	conv_row_47: 	reg_8bit port map (CLK => CLK, rst => '0', input => "110111100", output => elem_conv_row(47));
	conv_row_48: 	reg_8bit port map (CLK => CLK, rst => '0', input => "000111100", output => elem_conv_row(48));
	conv_row_49: 	reg_8bit port map (CLK => CLK, rst => '0', input => "001111100", output => elem_conv_row(49));
	conv_row_50: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111011111", output => elem_conv_row(50));
	conv_row_51: 	reg_8bit port map (CLK => CLK, rst => '0', input => "100001111", output => elem_conv_row(51));
	conv_row_52: 	reg_8bit port map (CLK => CLK, rst => '0', input => "100010111", output => elem_conv_row(52));
	conv_row_53: 	reg_8bit port map (CLK => CLK, rst => '0', input => "001110011", output => elem_conv_row(53));

	conv_row_54: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111100011", output => elem_conv_row(54));
	conv_row_55: 	reg_8bit port map (CLK => CLK, rst => '0', input => "101000011", output => elem_conv_row(55));
	conv_row_56: 	reg_8bit port map (CLK => CLK, rst => '0', input => "110001111", output => elem_conv_row(56));
	conv_row_57: 	reg_8bit port map (CLK => CLK, rst => '0', input => "100011111", output => elem_conv_row(57));
	conv_row_58: 	reg_8bit port map (CLK => CLK, rst => '0', input => "000111110", output => elem_conv_row(58));
	conv_row_59: 	reg_8bit port map (CLK => CLK, rst => '0', input => "001111110", output => elem_conv_row(59));
	conv_row_60: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111111100", output => elem_conv_row(60));
	conv_row_61: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111110011", output => elem_conv_row(61));
	conv_row_62: 	reg_8bit port map (CLK => CLK, rst => '0', input => "111000101", output => elem_conv_row(62));

	conv_row_63: 	reg_8bit port map (CLK => CLK, rst => '0', input => "010001100", output => elem_conv_row(63));
	conv_row_64: 	reg_8bit port map (CLK => CLK, rst => '0', input => "100011100", output => elem_conv_row(64));
	conv_row_65: 	reg_8bit port map (CLK => CLK, rst => '0', input => "001111010", output => elem_conv_row(65));
	conv_row_66: 	reg_8bit port map (CLK => CLK, rst => '0', input => "010011100", output => elem_conv_row(66));
	conv_row_67: 	reg_8bit port map (CLK => CLK, rst => '0', input => "000111000", output => elem_conv_row(67));
	conv_row_68: 	reg_8bit port map (CLK => CLK, rst => '0', input => "011111010", output => elem_conv_row(68));
	conv_row_69: 	reg_8bit port map (CLK => CLK, rst => '0', input => "000111000", output => elem_conv_row(69));
	conv_row_70: 	reg_8bit port map (CLK => CLK, rst => '0', input => "001111010", output => elem_conv_row(70));
	conv_row_71: 	reg_8bit port map (CLK => CLK, rst => '0', input => "010111100", output => elem_conv_row(71));

