	w_conv_0: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(0));
	w_conv_1: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(1));
	w_conv_2: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(2));
	w_conv_3: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(3));
	w_conv_4: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(4));
	w_conv_5: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(5));
	w_conv_6: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(6));
	w_conv_7: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(7));
	w_conv_8: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(8));
	w_conv_9: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(9));
	w_conv_10: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(10));
	w_conv_11: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(11));
	w_conv_12: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(12));
	w_conv_13: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(13));
	w_conv_14: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(14));
	w_conv_15: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(15));
	w_conv_16: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(16));
	w_conv_17: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(17));
	w_conv_18: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(18));
	w_conv_19: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(19));
	w_conv_20: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(20));
	w_conv_21: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(21));
	w_conv_22: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(22));
	w_conv_23: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(23));
	w_conv_24: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(24));
	w_conv_25: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(25));
	w_conv_26: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(26));
	w_conv_27: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(27));
	w_conv_28: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(28));
	w_conv_29: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(29));
	w_conv_30: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(30));
	w_conv_31: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(31));
	w_conv_32: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(32));
	w_conv_33: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(33));
	w_conv_34: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(34));
	w_conv_35: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(35));
	w_conv_36: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(36));
	w_conv_37: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(37));
	w_conv_38: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(38));
	w_conv_39: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(39));
	w_conv_40: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(40));
	w_conv_41: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(41));
	w_conv_42: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(42));
	w_conv_43: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(43));
	w_conv_44: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(44));
	w_conv_45: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(45));
	w_conv_46: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(46));
	w_conv_47: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(47));
	w_conv_48: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(48));
	w_conv_49: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(49));
	w_conv_50: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(50));
	w_conv_51: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(51));
	w_conv_52: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(52));
	w_conv_53: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(53));
	w_conv_54: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(54));
	w_conv_55: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(55));
	w_conv_56: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(56));
	w_conv_57: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(57));
	w_conv_58: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(58));
	w_conv_59: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(59));
	w_conv_60: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(60));
	w_conv_61: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(61));
	w_conv_62: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(62));
	w_conv_63: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(63));
	w_conv_64: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(64));
	w_conv_65: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(65));
	w_conv_66: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(66));
	w_conv_67: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(67));
	w_conv_68: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(68));
	w_conv_69: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(69));
	w_conv_70: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(70));
	w_conv_71: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(71));
	w_conv_72: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(72));
	w_conv_73: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(73));
	w_conv_74: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(74));
	w_conv_75: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(75));
	w_conv_76: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(76));
	w_conv_77: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(77));
	w_conv_78: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(78));
	w_conv_79: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(79));
	w_conv_80: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(80));

	w_conv_81: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(81));
	w_conv_82: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(82));
	w_conv_83: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(83));
	w_conv_84: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(84));
	w_conv_85: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(85));
	w_conv_86: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(86));
	w_conv_87: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(87));
	w_conv_88: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(88));
	w_conv_89: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(89));
	w_conv_90: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(90));
	w_conv_91: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(91));
	w_conv_92: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(92));
	w_conv_93: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(93));
	w_conv_94: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(94));
	w_conv_95: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(95));
	w_conv_96: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(96));
	w_conv_97: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(97));
	w_conv_98: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(98));
	w_conv_99: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(99));
	w_conv_100: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(100));
	w_conv_101: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(101));
	w_conv_102: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(102));
	w_conv_103: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(103));
	w_conv_104: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(104));
	w_conv_105: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(105));
	w_conv_106: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(106));
	w_conv_107: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(107));
	w_conv_108: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(108));
	w_conv_109: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(109));
	w_conv_110: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(110));
	w_conv_111: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(111));
	w_conv_112: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(112));
	w_conv_113: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(113));
	w_conv_114: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(114));
	w_conv_115: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(115));
	w_conv_116: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(116));
	w_conv_117: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(117));
	w_conv_118: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(118));
	w_conv_119: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(119));
	w_conv_120: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(120));
	w_conv_121: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(121));
	w_conv_122: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(122));
	w_conv_123: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(123));
	w_conv_124: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(124));
	w_conv_125: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(125));
	w_conv_126: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(126));
	w_conv_127: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(127));
	w_conv_128: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(128));
	w_conv_129: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(129));
	w_conv_130: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(130));
	w_conv_131: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(131));
	w_conv_132: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(132));
	w_conv_133: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(133));
	w_conv_134: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(134));
	w_conv_135: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(135));
	w_conv_136: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(136));
	w_conv_137: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(137));
	w_conv_138: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(138));
	w_conv_139: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(139));
	w_conv_140: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(140));
	w_conv_141: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(141));
	w_conv_142: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(142));
	w_conv_143: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(143));
	w_conv_144: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(144));
	w_conv_145: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(145));
	w_conv_146: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(146));
	w_conv_147: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(147));
	w_conv_148: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(148));
	w_conv_149: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(149));
	w_conv_150: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(150));
	w_conv_151: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(151));
	w_conv_152: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(152));
	w_conv_153: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(153));
	w_conv_154: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(154));
	w_conv_155: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(155));
	w_conv_156: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(156));
	w_conv_157: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(157));
	w_conv_158: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(158));
	w_conv_159: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(159));
	w_conv_160: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(160));
	w_conv_161: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(161));

	w_conv_162: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(162));
	w_conv_163: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(163));
	w_conv_164: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(164));
	w_conv_165: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(165));
	w_conv_166: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(166));
	w_conv_167: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(167));
	w_conv_168: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(168));
	w_conv_169: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(169));
	w_conv_170: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(170));
	w_conv_171: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(171));
	w_conv_172: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(172));
	w_conv_173: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(173));
	w_conv_174: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(174));
	w_conv_175: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(175));
	w_conv_176: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(176));
	w_conv_177: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(177));
	w_conv_178: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(178));
	w_conv_179: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(179));
	w_conv_180: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(180));
	w_conv_181: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(181));
	w_conv_182: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(182));
	w_conv_183: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(183));
	w_conv_184: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(184));
	w_conv_185: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(185));
	w_conv_186: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(186));
	w_conv_187: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(187));
	w_conv_188: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(188));
	w_conv_189: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(189));
	w_conv_190: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(190));
	w_conv_191: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(191));
	w_conv_192: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(192));
	w_conv_193: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(193));
	w_conv_194: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(194));
	w_conv_195: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(195));
	w_conv_196: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(196));
	w_conv_197: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(197));
	w_conv_198: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(198));
	w_conv_199: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(199));
	w_conv_200: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(200));
	w_conv_201: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(201));
	w_conv_202: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(202));
	w_conv_203: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(203));
	w_conv_204: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(204));
	w_conv_205: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(205));
	w_conv_206: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(206));
	w_conv_207: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(207));
	w_conv_208: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(208));
	w_conv_209: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(209));
	w_conv_210: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(210));
	w_conv_211: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(211));
	w_conv_212: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(212));
	w_conv_213: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(213));
	w_conv_214: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(214));
	w_conv_215: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(215));
	w_conv_216: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(216));
	w_conv_217: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(217));
	w_conv_218: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(218));
	w_conv_219: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(219));
	w_conv_220: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(220));
	w_conv_221: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(221));
	w_conv_222: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(222));
	w_conv_223: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(223));
	w_conv_224: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(224));
	w_conv_225: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(225));
	w_conv_226: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(226));
	w_conv_227: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(227));
	w_conv_228: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(228));
	w_conv_229: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(229));
	w_conv_230: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(230));
	w_conv_231: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(231));
	w_conv_232: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(232));
	w_conv_233: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(233));
	w_conv_234: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(234));
	w_conv_235: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(235));
	w_conv_236: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(236));
	w_conv_237: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(237));
	w_conv_238: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(238));
	w_conv_239: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(239));
	w_conv_240: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(240));
	w_conv_241: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(241));
	w_conv_242: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(242));

	w_conv_243: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(243));
	w_conv_244: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(244));
	w_conv_245: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(245));
	w_conv_246: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(246));
	w_conv_247: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(247));
	w_conv_248: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(248));
	w_conv_249: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(249));
	w_conv_250: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(250));
	w_conv_251: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(251));
	w_conv_252: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(252));
	w_conv_253: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(253));
	w_conv_254: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(254));
	w_conv_255: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(255));
	w_conv_256: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(256));
	w_conv_257: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(257));
	w_conv_258: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(258));
	w_conv_259: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(259));
	w_conv_260: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(260));
	w_conv_261: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(261));
	w_conv_262: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(262));
	w_conv_263: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(263));
	w_conv_264: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(264));
	w_conv_265: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(265));
	w_conv_266: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(266));
	w_conv_267: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(267));
	w_conv_268: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(268));
	w_conv_269: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(269));
	w_conv_270: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(270));
	w_conv_271: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(271));
	w_conv_272: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(272));
	w_conv_273: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(273));
	w_conv_274: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(274));
	w_conv_275: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(275));
	w_conv_276: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(276));
	w_conv_277: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(277));
	w_conv_278: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(278));
	w_conv_279: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(279));
	w_conv_280: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(280));
	w_conv_281: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(281));
	w_conv_282: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(282));
	w_conv_283: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(283));
	w_conv_284: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(284));
	w_conv_285: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(285));
	w_conv_286: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(286));
	w_conv_287: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(287));
	w_conv_288: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(288));
	w_conv_289: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(289));
	w_conv_290: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(290));
	w_conv_291: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(291));
	w_conv_292: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(292));
	w_conv_293: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(293));
	w_conv_294: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(294));
	w_conv_295: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(295));
	w_conv_296: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(296));
	w_conv_297: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(297));
	w_conv_298: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(298));
	w_conv_299: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(299));
	w_conv_300: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(300));
	w_conv_301: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(301));
	w_conv_302: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(302));
	w_conv_303: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(303));
	w_conv_304: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(304));
	w_conv_305: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(305));
	w_conv_306: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(306));
	w_conv_307: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(307));
	w_conv_308: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(308));
	w_conv_309: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(309));
	w_conv_310: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(310));
	w_conv_311: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(311));
	w_conv_312: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(312));
	w_conv_313: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(313));
	w_conv_314: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(314));
	w_conv_315: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(315));
	w_conv_316: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(316));
	w_conv_317: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(317));
	w_conv_318: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(318));
	w_conv_319: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(319));
	w_conv_320: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(320));
	w_conv_321: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(321));
	w_conv_322: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(322));
	w_conv_323: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(323));

	w_conv_324: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(324));
	w_conv_325: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(325));
	w_conv_326: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(326));
	w_conv_327: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(327));
	w_conv_328: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(328));
	w_conv_329: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(329));
	w_conv_330: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(330));
	w_conv_331: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(331));
	w_conv_332: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(332));
	w_conv_333: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(333));
	w_conv_334: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(334));
	w_conv_335: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(335));
	w_conv_336: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(336));
	w_conv_337: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(337));
	w_conv_338: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(338));
	w_conv_339: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(339));
	w_conv_340: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(340));
	w_conv_341: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(341));
	w_conv_342: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(342));
	w_conv_343: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(343));
	w_conv_344: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(344));
	w_conv_345: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(345));
	w_conv_346: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(346));
	w_conv_347: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(347));
	w_conv_348: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(348));
	w_conv_349: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(349));
	w_conv_350: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(350));
	w_conv_351: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(351));
	w_conv_352: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(352));
	w_conv_353: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(353));
	w_conv_354: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(354));
	w_conv_355: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(355));
	w_conv_356: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(356));
	w_conv_357: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(357));
	w_conv_358: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(358));
	w_conv_359: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(359));
	w_conv_360: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(360));
	w_conv_361: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(361));
	w_conv_362: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(362));
	w_conv_363: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(363));
	w_conv_364: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(364));
	w_conv_365: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(365));
	w_conv_366: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(366));
	w_conv_367: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(367));
	w_conv_368: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(368));
	w_conv_369: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(369));
	w_conv_370: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(370));
	w_conv_371: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(371));
	w_conv_372: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(372));
	w_conv_373: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(373));
	w_conv_374: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(374));
	w_conv_375: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(375));
	w_conv_376: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(376));
	w_conv_377: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(377));
	w_conv_378: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(378));
	w_conv_379: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(379));
	w_conv_380: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(380));
	w_conv_381: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(381));
	w_conv_382: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(382));
	w_conv_383: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(383));
	w_conv_384: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(384));
	w_conv_385: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(385));
	w_conv_386: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(386));
	w_conv_387: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(387));
	w_conv_388: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(388));
	w_conv_389: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(389));
	w_conv_390: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(390));
	w_conv_391: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(391));
	w_conv_392: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(392));
	w_conv_393: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(393));
	w_conv_394: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(394));
	w_conv_395: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(395));
	w_conv_396: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(396));
	w_conv_397: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(397));
	w_conv_398: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(398));
	w_conv_399: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(399));
	w_conv_400: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(400));
	w_conv_401: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(401));
	w_conv_402: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(402));
	w_conv_403: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(403));
	w_conv_404: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(404));

	w_conv_405: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(405));
	w_conv_406: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(406));
	w_conv_407: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(407));
	w_conv_408: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(408));
	w_conv_409: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(409));
	w_conv_410: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(410));
	w_conv_411: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(411));
	w_conv_412: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(412));
	w_conv_413: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(413));
	w_conv_414: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(414));
	w_conv_415: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(415));
	w_conv_416: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(416));
	w_conv_417: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(417));
	w_conv_418: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(418));
	w_conv_419: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(419));
	w_conv_420: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(420));
	w_conv_421: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(421));
	w_conv_422: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(422));
	w_conv_423: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(423));
	w_conv_424: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(424));
	w_conv_425: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(425));
	w_conv_426: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(426));
	w_conv_427: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(427));
	w_conv_428: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(428));
	w_conv_429: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(429));
	w_conv_430: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(430));
	w_conv_431: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(431));
	w_conv_432: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(432));
	w_conv_433: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(433));
	w_conv_434: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(434));
	w_conv_435: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(435));
	w_conv_436: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(436));
	w_conv_437: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(437));
	w_conv_438: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(438));
	w_conv_439: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(439));
	w_conv_440: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(440));
	w_conv_441: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(441));
	w_conv_442: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(442));
	w_conv_443: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(443));
	w_conv_444: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(444));
	w_conv_445: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(445));
	w_conv_446: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(446));
	w_conv_447: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(447));
	w_conv_448: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(448));
	w_conv_449: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(449));
	w_conv_450: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(450));
	w_conv_451: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(451));
	w_conv_452: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(452));
	w_conv_453: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(453));
	w_conv_454: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(454));
	w_conv_455: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(455));
	w_conv_456: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(456));
	w_conv_457: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(457));
	w_conv_458: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(458));
	w_conv_459: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(459));
	w_conv_460: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(460));
	w_conv_461: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(461));
	w_conv_462: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(462));
	w_conv_463: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(463));
	w_conv_464: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(464));
	w_conv_465: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(465));
	w_conv_466: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(466));
	w_conv_467: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(467));
	w_conv_468: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(468));
	w_conv_469: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(469));
	w_conv_470: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(470));
	w_conv_471: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(471));
	w_conv_472: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(472));
	w_conv_473: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(473));
	w_conv_474: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(474));
	w_conv_475: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(475));
	w_conv_476: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(476));
	w_conv_477: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(477));
	w_conv_478: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(478));
	w_conv_479: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(479));
	w_conv_480: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(480));
	w_conv_481: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(481));
	w_conv_482: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(482));
	w_conv_483: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(483));
	w_conv_484: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(484));
	w_conv_485: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(485));

	w_conv_486: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(486));
	w_conv_487: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(487));
	w_conv_488: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(488));
	w_conv_489: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(489));
	w_conv_490: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(490));
	w_conv_491: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(491));
	w_conv_492: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(492));
	w_conv_493: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(493));
	w_conv_494: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(494));
	w_conv_495: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(495));
	w_conv_496: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(496));
	w_conv_497: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(497));
	w_conv_498: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(498));
	w_conv_499: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(499));
	w_conv_500: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(500));
	w_conv_501: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(501));
	w_conv_502: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(502));
	w_conv_503: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(503));
	w_conv_504: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(504));
	w_conv_505: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(505));
	w_conv_506: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(506));
	w_conv_507: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(507));
	w_conv_508: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(508));
	w_conv_509: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(509));
	w_conv_510: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(510));
	w_conv_511: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(511));
	w_conv_512: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(512));
	w_conv_513: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(513));
	w_conv_514: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(514));
	w_conv_515: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(515));
	w_conv_516: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(516));
	w_conv_517: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(517));
	w_conv_518: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(518));
	w_conv_519: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(519));
	w_conv_520: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(520));
	w_conv_521: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(521));
	w_conv_522: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(522));
	w_conv_523: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(523));
	w_conv_524: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(524));
	w_conv_525: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(525));
	w_conv_526: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(526));
	w_conv_527: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(527));
	w_conv_528: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(528));
	w_conv_529: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(529));
	w_conv_530: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(530));
	w_conv_531: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(531));
	w_conv_532: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(532));
	w_conv_533: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(533));
	w_conv_534: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(534));
	w_conv_535: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(535));
	w_conv_536: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(536));
	w_conv_537: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(537));
	w_conv_538: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(538));
	w_conv_539: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(539));
	w_conv_540: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(540));
	w_conv_541: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(541));
	w_conv_542: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(542));
	w_conv_543: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(543));
	w_conv_544: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(544));
	w_conv_545: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(545));
	w_conv_546: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(546));
	w_conv_547: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(547));
	w_conv_548: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(548));
	w_conv_549: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(549));
	w_conv_550: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(550));
	w_conv_551: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(551));
	w_conv_552: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(552));
	w_conv_553: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(553));
	w_conv_554: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(554));
	w_conv_555: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(555));
	w_conv_556: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(556));
	w_conv_557: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(557));
	w_conv_558: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(558));
	w_conv_559: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(559));
	w_conv_560: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(560));
	w_conv_561: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(561));
	w_conv_562: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(562));
	w_conv_563: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(563));
	w_conv_564: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(564));
	w_conv_565: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(565));
	w_conv_566: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(566));

	w_conv_567: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(567));
	w_conv_568: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(568));
	w_conv_569: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(569));
	w_conv_570: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(570));
	w_conv_571: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(571));
	w_conv_572: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(572));
	w_conv_573: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(573));
	w_conv_574: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(574));
	w_conv_575: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(575));
	w_conv_576: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(576));
	w_conv_577: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(577));
	w_conv_578: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(578));
	w_conv_579: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(579));
	w_conv_580: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(580));
	w_conv_581: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(581));
	w_conv_582: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(582));
	w_conv_583: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(583));
	w_conv_584: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(584));
	w_conv_585: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(585));
	w_conv_586: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(586));
	w_conv_587: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(587));
	w_conv_588: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(588));
	w_conv_589: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(589));
	w_conv_590: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(590));
	w_conv_591: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(591));
	w_conv_592: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(592));
	w_conv_593: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(593));
	w_conv_594: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(594));
	w_conv_595: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(595));
	w_conv_596: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(596));
	w_conv_597: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(597));
	w_conv_598: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(598));
	w_conv_599: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(599));
	w_conv_600: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(600));
	w_conv_601: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(601));
	w_conv_602: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(602));
	w_conv_603: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(603));
	w_conv_604: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(604));
	w_conv_605: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(605));
	w_conv_606: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(606));
	w_conv_607: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(607));
	w_conv_608: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(608));
	w_conv_609: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(609));
	w_conv_610: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(610));
	w_conv_611: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(611));
	w_conv_612: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(612));
	w_conv_613: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(613));
	w_conv_614: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(614));
	w_conv_615: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(615));
	w_conv_616: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(616));
	w_conv_617: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(617));
	w_conv_618: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(618));
	w_conv_619: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(619));
	w_conv_620: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(620));
	w_conv_621: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(621));
	w_conv_622: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(622));
	w_conv_623: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(623));
	w_conv_624: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(624));
	w_conv_625: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(625));
	w_conv_626: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(626));
	w_conv_627: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(627));
	w_conv_628: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(628));
	w_conv_629: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(629));
	w_conv_630: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(630));
	w_conv_631: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(631));
	w_conv_632: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(632));
	w_conv_633: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(633));
	w_conv_634: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(634));
	w_conv_635: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(635));
	w_conv_636: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(636));
	w_conv_637: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(637));
	w_conv_638: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(638));
	w_conv_639: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(639));
	w_conv_640: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(640));
	w_conv_641: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(641));
	w_conv_642: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(642));
	w_conv_643: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(643));
	w_conv_644: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(644));
	w_conv_645: 	reg_8bit port map (CLK => CLK, rst => '0', input => '1', output => elem_w_conv(645));
	w_conv_646: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(646));
	w_conv_647: 	reg_8bit port map (CLK => CLK, rst => '0', input => '0', output => elem_w_conv(647));

