	img_row_0: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000000000000000000000", output => elem_img_row(0));
	img_row_1: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000000000000000000000", output => elem_img_row(1));
	img_row_2: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000000000000000000000", output => elem_img_row(2));
	img_row_3: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000000000000000000000", output => elem_img_row(3));
	img_row_4: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000001111100000000000", output => elem_img_row(4));
	img_row_5: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000111111110000000000", output => elem_img_row(5));
	img_row_6: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000001111111110000000000", output => elem_img_row(6));
	img_row_7: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000000001110000000000", output => elem_img_row(7));
	img_row_8: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000000011110000000000", output => elem_img_row(8));
	img_row_9: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000000011100000000000", output => elem_img_row(9));
	img_row_10: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000000111000000000000", output => elem_img_row(10));
	img_row_11: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000001110000000000000", output => elem_img_row(11));
	img_row_12: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000011111000000000000", output => elem_img_row(12));
	img_row_13: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000011111100000000000", output => elem_img_row(13));
	img_row_14: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000000111110000000000", output => elem_img_row(14));
	img_row_15: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000000001111000000000", output => elem_img_row(15));
	img_row_16: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000000000111000000000", output => elem_img_row(16));
	img_row_17: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000000000011100000000", output => elem_img_row(17));
	img_row_18: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000000000011100000000", output => elem_img_row(18));
	img_row_19: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000000000011100000000", output => elem_img_row(19));
	img_row_20: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000011000001111000000000", output => elem_img_row(20));
	img_row_21: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000011111111110000000000", output => elem_img_row(21));
	img_row_22: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000011111111100000000000", output => elem_img_row(22));
	img_row_23: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000111000000000000000", output => elem_img_row(23));
	img_row_24: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000000000000000000000", output => elem_img_row(24));
	img_row_25: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000000000000000000000", output => elem_img_row(25));
	img_row_26: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000000000000000000000", output => elem_img_row(26));
	img_row_27: 	reg_8bit port map (CLK => CLK, rst => '0', input => "0000000000000000000000000000", output => elem_img_row(27));
